interface uart_rx_intf();
    logic clk;
    logic reset_n;
    logic rts_n;
    logic rx;
endinterface