
`define DATA_5BIT 2'b00
`define DATA_6BIT 2'b01
`define DATA_7BIT 2'b10
`define DATA_8BIT 2'b11
typedef logic [ 7 : 0] uart