interface uart_tx_intf();
    logic clk;
    logic reset_n;
    logic cts_n;
    logic tx;
endinterface