class uart_rx_transaction extends uvm_object