`include "uvm.sv"
`include "uvm_macros.svh"
import uvm_pkg::*;

//`include "uart_env"
`include "define.sv"
`include "uart_sw_intf.sv"
`include "uart_sw_item.sv"
`include "uart_sw_sequencer.sv"
`include "uart_sequence.sv"
`include "uart_standard_send_seq.sv"
`include "uart_sw_monitor.sv"
`include "uart_sw_driver.sv"
`include "uart_sw_agent.sv"
// `include "dti_uart_env.sv"

// `include "dti_uart_tx_seq.sv"
// `include "dti_uart_rx_seq.sv"

// `include "dti_uart_base_test.sv"
// `include "dti_uart_random_test.sv"