//include UVM
`include "uvm.sv"
`include "uvm_macros.svh"
import uvm_pkg::*;
//include Package
`include "include_files.sv"

//include environment
`include "uart_env.sv"

//include sequence apb


//include sequence uart

//include test
`include "uart_test.sv"

