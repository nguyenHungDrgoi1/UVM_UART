
`define DATA_5BIT 2'b00
`define DATA_6BIT 2'b01
`define DATA_7BIT 2'b10
`define DATA_8BIT 2'b11
`define DATA_FRAME_5BIT 5
`define DATA_FRAME_6BIT 6
`define DATA_FRAME_7BIT 7
`define DATA_FRAME_8BIT 8
`define UART_PARITY_ODD 0
`define UART_TWO_STOP_BIT 1
typedef logic [ 7 : 0] uart_data_frame;
//fill note